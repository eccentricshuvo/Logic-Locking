// Benchmark "s1196_xor" written by ABC on Thu Oct 21 13:39:17 2021

module s1196_xor ( clock, 
    G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, keyinput0,
    keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
    keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
    keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
    keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
    keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30,
    keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36,
    keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
    keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
    keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
    keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60,
    keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66,
    keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
    keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
    keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
    keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90,
    keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96,
    keyinput97, keyinput98, keyinput99, keyinput100, keyinput101,
    keyinput102, keyinput103, keyinput104, keyinput105, keyinput106,
    keyinput107, keyinput108, keyinput109, keyinput110, keyinput111,
    keyinput112, keyinput113, keyinput114, keyinput115, keyinput116,
    keyinput117, keyinput118, keyinput119, keyinput120, keyinput121,
    keyinput122, keyinput123, keyinput124, keyinput125, keyinput126,
    keyinput127,
    G546, G539, G550, G551, G552, G547, G548, G549, G530, G45, G542, G532,
    G535, G537  );
  input  clock;
  input  G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13,
    keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5,
    keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11,
    keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
    keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
    keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
    keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35,
    keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41,
    keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
    keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
    keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
    keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65,
    keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71,
    keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
    keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
    keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
    keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95,
    keyinput96, keyinput97, keyinput98, keyinput99, keyinput100,
    keyinput101, keyinput102, keyinput103, keyinput104, keyinput105,
    keyinput106, keyinput107, keyinput108, keyinput109, keyinput110,
    keyinput111, keyinput112, keyinput113, keyinput114, keyinput115,
    keyinput116, keyinput117, keyinput118, keyinput119, keyinput120,
    keyinput121, keyinput122, keyinput123, keyinput124, keyinput125,
    keyinput126, keyinput127;
  output G546, G539, G550, G551, G552, G547, G548, G549, G530, G45, G542,
    G532, G535, G537;
  reg G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46;
  wire new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_1_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_1_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_1_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_1_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_1_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_1_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_1_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_1_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_1_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_1_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_1_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_1_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_1_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_1_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_1_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_1_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_1_, new_n395_, new_n396_,
    new_n397_, new_n398_1_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n955_, new_n956_, new_n957_, new_n958_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n976_, new_n979_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, n314, n319, n324, n329,
    n334, n339, n344, n349, n354, n359, n364, n369, n374, n379, n384, n389,
    n394, n398;
  assign new_n211_ = ~G7 & G8;
  assign new_n212_ = keyinput23 & new_n211_;
  assign new_n213_ = ~keyinput23 & ~new_n211_;
  assign new_n214_ = ~new_n212_ & ~new_n213_;
  assign new_n215_ = ~G10 & keyinput0;
  assign new_n216_ = G10 & ~keyinput0;
  assign new_n217_ = ~new_n215_ & ~new_n216_;
  assign new_n218_ = G9 & ~new_n217_;
  assign new_n219_ = ~new_n214_ & new_n218_;
  assign new_n220_ = keyinput22 & ~new_n219_;
  assign new_n221_ = ~keyinput22 & new_n219_;
  assign new_n222_ = ~new_n220_ & ~new_n221_;
  assign new_n223_ = ~G8 & G10;
  assign new_n224_ = ~G7 & G9;
  assign new_n225_ = new_n223_ & new_n224_;
  assign new_n226_ = G7 & ~G10;
  assign new_n227_ = ~G9 & new_n226_;
  assign new_n228_ = G8 & new_n227_;
  assign new_n229_ = ~new_n225_ & ~new_n228_;
  assign new_n230_ = new_n222_ & new_n229_;
  assign new_n231_ = ~G11 & keyinput12;
  assign new_n232_ = G11 & ~keyinput12;
  assign new_n233_ = ~new_n231_ & ~new_n232_;
  assign new_n234_ = G4 & G6;
  assign new_n235_ = G3 & new_n234_;
  assign new_n236_ = ~G5 & new_n233_;
  assign new_n237_ = new_n235_ & new_n236_;
  assign new_n238_ = keyinput7 & ~new_n237_;
  assign new_n239_ = ~keyinput7 & new_n237_;
  assign new_n240_ = ~new_n238_ & ~new_n239_;
  assign new_n241_ = ~G2 & ~new_n230_;
  assign new_n242_ = ~new_n240_ & new_n241_;
  assign new_n243_ = G3 & G5;
  assign new_n244_ = G9 & G11;
  assign new_n245_ = keyinput53 & ~new_n244_;
  assign new_n246_ = ~keyinput53 & new_n244_;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign new_n248_ = G8 & ~new_n247_;
  assign new_n249_ = G7 & G10;
  assign new_n250_ = new_n248_ & new_n249_;
  assign new_n251_ = new_n234_ & new_n243_;
  assign new_n252_ = new_n250_ & new_n251_;
  assign new_n253_ = ~G4 & ~G5;
  assign new_n254_ = G3 & G11;
  assign new_n255_ = G35 & new_n254_;
  assign new_n256_ = new_n253_ & new_n255_;
  assign new_n257_ = keyinput103 & ~new_n256_;
  assign new_n258_ = ~keyinput103 & new_n256_;
  assign new_n259_ = ~new_n257_ & ~new_n258_;
  assign new_n260_ = ~G7 & ~G11;
  assign new_n261_ = ~G8 & new_n260_;
  assign new_n262_ = keyinput121 & new_n261_;
  assign new_n263_ = ~keyinput121 & ~new_n261_;
  assign new_n264_ = ~new_n262_ & ~new_n263_;
  assign new_n265_ = new_n218_ & ~new_n264_;
  assign new_n266_ = G5 & new_n265_;
  assign new_n267_ = new_n235_ & new_n266_;
  assign new_n268_ = ~new_n252_ & ~new_n259_;
  assign new_n269_ = ~new_n267_ & new_n268_;
  assign new_n270_ = keyinput34 & ~new_n269_;
  assign new_n271_ = ~keyinput34 & new_n269_;
  assign new_n272_ = ~new_n270_ & ~new_n271_;
  assign new_n273_ = G2 & ~new_n272_;
  assign new_n274_ = keyinput57 & ~new_n273_;
  assign new_n275_ = ~keyinput57 & new_n273_;
  assign new_n276_ = ~new_n274_ & ~new_n275_;
  assign new_n277_ = ~G6 & G36;
  assign new_n278_ = G5 & new_n234_;
  assign new_n279_ = keyinput5 & new_n278_;
  assign new_n280_ = ~keyinput5 & ~new_n278_;
  assign new_n281_ = ~new_n279_ & ~new_n280_;
  assign new_n282_ = G11 & ~new_n229_;
  assign new_n283_ = ~new_n281_ & new_n282_;
  assign new_n284_ = ~new_n277_ & ~new_n283_;
  assign new_n285_ = ~G3 & ~new_n284_;
  assign new_n286_ = keyinput115 & new_n285_;
  assign new_n287_ = ~keyinput115 & ~new_n285_;
  assign new_n288_ = ~new_n286_ & ~new_n287_;
  assign new_n289_ = ~G2 & ~new_n288_;
  assign new_n290_ = ~new_n242_ & new_n276_;
  assign new_n291_ = ~new_n289_ & new_n290_;
  assign new_n292_ = G30 & new_n211_;
  assign new_n293_ = ~new_n248_ & new_n249_;
  assign new_n294_ = G7 & new_n218_;
  assign new_n295_ = ~new_n292_ & ~new_n293_;
  assign new_n296_ = ~new_n294_ & new_n295_;
  assign new_n297_ = keyinput47 & G32;
  assign new_n298_ = ~keyinput47 & ~G32;
  assign new_n299_ = ~new_n297_ & ~new_n298_;
  assign new_n300_ = ~new_n296_ & ~new_n299_;
  assign new_n301_ = keyinput27 & ~new_n300_;
  assign new_n302_ = ~keyinput27 & new_n300_;
  assign new_n303_ = ~new_n301_ & ~new_n302_;
  assign new_n304_ = keyinput82 & new_n303_;
  assign new_n305_ = ~keyinput82 & ~new_n303_;
  assign new_n306_ = ~new_n304_ & ~new_n305_;
  assign new_n307_ = ~G13 & new_n306_;
  assign new_n308_ = ~G12 & new_n291_;
  assign new_n309_ = new_n307_ & new_n308_;
  assign new_n310_ = keyinput105 & ~new_n309_;
  assign new_n311_ = ~keyinput105 & new_n309_;
  assign new_n312_ = ~new_n310_ & ~new_n311_;
  assign new_n313_ = ~G5 & ~G7;
  assign new_n314_1_ = keyinput91 & ~new_n223_;
  assign new_n315_ = ~keyinput91 & new_n223_;
  assign new_n316_ = ~new_n314_1_ & ~new_n315_;
  assign new_n317_ = G6 & ~G9;
  assign new_n318_ = ~G3 & new_n313_;
  assign new_n319_1_ = ~new_n316_ & new_n318_;
  assign new_n320_ = new_n317_ & new_n319_1_;
  assign new_n321_ = G8 & new_n243_;
  assign new_n322_ = G37 & new_n321_;
  assign new_n323_ = new_n226_ & new_n322_;
  assign new_n324_1_ = ~new_n320_ & ~new_n323_;
  assign new_n325_ = keyinput113 & new_n324_1_;
  assign new_n326_ = ~keyinput113 & ~new_n324_1_;
  assign new_n327_ = ~new_n325_ & ~new_n326_;
  assign new_n328_ = ~G0 & ~G4;
  assign new_n329_1_ = G11 & ~new_n327_;
  assign new_n330_ = new_n328_ & new_n329_1_;
  assign new_n331_ = keyinput16 & ~new_n330_;
  assign new_n332_ = ~keyinput16 & new_n330_;
  assign new_n333_ = ~new_n331_ & ~new_n332_;
  assign new_n334_1_ = G0 & new_n252_;
  assign new_n335_ = new_n333_ & ~new_n334_1_;
  assign new_n336_ = G1 & G2;
  assign new_n337_ = ~new_n335_ & new_n336_;
  assign new_n338_ = keyinput13 & new_n337_;
  assign new_n339_1_ = ~keyinput13 & ~new_n337_;
  assign new_n340_ = ~new_n338_ & ~new_n339_1_;
  assign new_n341_ = keyinput50 & G46;
  assign new_n342_ = ~keyinput50 & ~G46;
  assign new_n343_ = ~new_n341_ & ~new_n342_;
  assign new_n344_1_ = ~G10 & ~G11;
  assign new_n345_ = keyinput48 & new_n344_1_;
  assign new_n346_ = ~keyinput48 & ~new_n344_1_;
  assign new_n347_ = ~new_n345_ & ~new_n346_;
  assign new_n348_ = ~G9 & new_n347_;
  assign new_n349_1_ = ~G6 & G7;
  assign new_n350_ = G30 & new_n349_1_;
  assign new_n351_ = G8 & G31;
  assign new_n352_ = keyinput112 & ~new_n351_;
  assign new_n353_ = ~keyinput112 & new_n351_;
  assign new_n354_1_ = ~new_n352_ & ~new_n353_;
  assign new_n355_ = new_n348_ & ~new_n350_;
  assign new_n356_ = ~new_n354_1_ & new_n355_;
  assign new_n357_ = keyinput54 & new_n356_;
  assign new_n358_ = ~keyinput54 & ~new_n356_;
  assign new_n359_1_ = ~new_n357_ & ~new_n358_;
  assign new_n360_ = G8 & ~G31;
  assign new_n361_ = ~new_n223_ & ~new_n360_;
  assign new_n362_ = G9 & ~new_n361_;
  assign new_n363_ = new_n260_ & new_n362_;
  assign new_n364_1_ = keyinput56 & ~new_n363_;
  assign new_n365_ = ~keyinput56 & new_n363_;
  assign new_n366_ = ~new_n364_1_ & ~new_n365_;
  assign new_n367_ = G8 & G10;
  assign new_n368_ = G9 & ~new_n367_;
  assign new_n369_1_ = keyinput111 & new_n360_;
  assign new_n370_ = ~keyinput111 & ~new_n360_;
  assign new_n371_ = ~new_n369_1_ & ~new_n370_;
  assign new_n372_ = ~new_n350_ & ~new_n368_;
  assign new_n373_ = ~new_n371_ & new_n372_;
  assign new_n374_1_ = ~G6 & ~G30;
  assign new_n375_ = ~G7 & ~G8;
  assign new_n376_ = keyinput127 & new_n375_;
  assign new_n377_ = ~keyinput127 & ~new_n375_;
  assign new_n378_ = ~new_n376_ & ~new_n377_;
  assign new_n379_1_ = ~G9 & ~new_n378_;
  assign new_n380_ = ~new_n373_ & ~new_n374_1_;
  assign new_n381_ = ~new_n379_1_ & new_n380_;
  assign new_n382_ = G11 & ~new_n381_;
  assign new_n383_ = G3 & new_n328_;
  assign new_n384_1_ = ~G1 & G5;
  assign new_n385_ = G4 & ~new_n243_;
  assign new_n386_ = ~new_n384_1_ & ~new_n385_;
  assign new_n387_ = keyinput96 & new_n386_;
  assign new_n388_ = ~keyinput96 & ~new_n386_;
  assign new_n389_1_ = ~new_n387_ & ~new_n388_;
  assign new_n390_ = G2 & new_n389_1_;
  assign new_n391_ = ~G3 & ~new_n390_;
  assign new_n392_ = keyinput120 & ~new_n391_;
  assign new_n393_ = ~keyinput120 & new_n391_;
  assign new_n394_1_ = ~new_n392_ & ~new_n393_;
  assign new_n395_ = ~G5 & new_n394_1_;
  assign new_n396_ = ~new_n383_ & ~new_n395_;
  assign new_n397_ = G4 & ~G5;
  assign new_n398_1_ = ~new_n396_ & ~new_n397_;
  assign new_n399_ = keyinput49 & ~new_n398_1_;
  assign new_n400_ = ~keyinput49 & new_n398_1_;
  assign new_n401_ = ~new_n399_ & ~new_n400_;
  assign new_n402_ = new_n359_1_ & new_n366_;
  assign new_n403_ = ~new_n382_ & new_n402_;
  assign new_n404_ = new_n401_ & new_n403_;
  assign new_n405_ = keyinput55 & ~new_n404_;
  assign new_n406_ = ~keyinput55 & new_n404_;
  assign new_n407_ = ~new_n405_ & ~new_n406_;
  assign new_n408_ = ~new_n343_ & ~new_n407_;
  assign new_n409_ = keyinput97 & ~new_n408_;
  assign new_n410_ = ~keyinput97 & new_n408_;
  assign new_n411_ = ~new_n409_ & ~new_n410_;
  assign new_n412_ = G12 & ~G13;
  assign new_n413_ = ~new_n411_ & new_n412_;
  assign new_n414_ = keyinput118 & new_n413_;
  assign new_n415_ = ~keyinput118 & ~new_n413_;
  assign new_n416_ = ~new_n414_ & ~new_n415_;
  assign new_n417_ = ~new_n340_ & ~new_n416_;
  assign new_n418_ = keyinput81 & ~new_n417_;
  assign new_n419_ = ~keyinput81 & new_n417_;
  assign new_n420_ = ~new_n418_ & ~new_n419_;
  assign new_n421_ = G1 & G3;
  assign new_n422_ = ~G4 & new_n421_;
  assign new_n423_ = G6 & new_n422_;
  assign new_n424_ = ~G1 & new_n235_;
  assign new_n425_ = ~new_n423_ & ~new_n424_;
  assign new_n426_ = ~new_n247_ & ~new_n316_;
  assign new_n427_ = keyinput68 & ~new_n426_;
  assign new_n428_ = ~keyinput68 & new_n426_;
  assign new_n429_ = ~new_n427_ & ~new_n428_;
  assign new_n430_ = keyinput95 & new_n429_;
  assign new_n431_ = ~keyinput95 & ~new_n429_;
  assign new_n432_ = ~new_n430_ & ~new_n431_;
  assign new_n433_ = ~new_n425_ & ~new_n432_;
  assign new_n434_ = ~G10 & new_n248_;
  assign new_n435_ = keyinput83 & ~new_n434_;
  assign new_n436_ = ~keyinput83 & new_n434_;
  assign new_n437_ = ~new_n435_ & ~new_n436_;
  assign new_n438_ = new_n424_ & ~new_n437_;
  assign new_n439_ = ~new_n433_ & ~new_n438_;
  assign new_n440_ = ~G7 & ~new_n439_;
  assign new_n441_ = ~G4 & ~G6;
  assign new_n442_ = ~G1 & G3;
  assign new_n443_ = ~G8 & new_n441_;
  assign new_n444_ = new_n442_ & new_n443_;
  assign new_n445_ = G8 & ~new_n425_;
  assign new_n446_ = ~new_n444_ & ~new_n445_;
  assign new_n447_ = new_n227_ & new_n233_;
  assign new_n448_ = ~new_n446_ & new_n447_;
  assign new_n449_ = ~new_n440_ & ~new_n448_;
  assign new_n450_ = G2 & ~G5;
  assign new_n451_ = ~new_n449_ & new_n450_;
  assign new_n452_ = ~new_n250_ & ~new_n265_;
  assign new_n453_ = G2 & new_n234_;
  assign new_n454_ = G1 & new_n243_;
  assign new_n455_ = ~new_n452_ & new_n453_;
  assign new_n456_ = new_n454_ & new_n455_;
  assign new_n457_ = keyinput19 & ~new_n456_;
  assign new_n458_ = ~keyinput19 & new_n456_;
  assign new_n459_ = ~new_n457_ & ~new_n458_;
  assign new_n460_ = ~new_n451_ & new_n459_;
  assign new_n461_ = ~G3 & new_n397_;
  assign new_n462_ = keyinput4 & ~new_n461_;
  assign new_n463_ = ~keyinput4 & new_n461_;
  assign new_n464_ = ~new_n462_ & ~new_n463_;
  assign new_n465_ = ~G2 & G3;
  assign new_n466_ = G2 & ~G3;
  assign new_n467_ = ~new_n465_ & ~new_n466_;
  assign new_n468_ = ~new_n385_ & new_n467_;
  assign new_n469_ = G6 & ~new_n468_;
  assign new_n470_ = keyinput99 & new_n469_;
  assign new_n471_ = ~keyinput99 & ~new_n469_;
  assign new_n472_ = ~new_n470_ & ~new_n471_;
  assign new_n473_ = G3 & ~new_n234_;
  assign new_n474_ = ~new_n441_ & ~new_n473_;
  assign new_n475_ = G5 & ~new_n474_;
  assign new_n476_ = new_n464_ & new_n472_;
  assign new_n477_ = ~new_n475_ & new_n476_;
  assign new_n478_ = G1 & ~new_n477_;
  assign new_n479_ = G1 & G4;
  assign new_n480_ = keyinput109 & ~new_n479_;
  assign new_n481_ = ~keyinput109 & new_n479_;
  assign new_n482_ = ~new_n480_ & ~new_n481_;
  assign new_n483_ = G2 & new_n482_;
  assign new_n484_ = ~G6 & new_n483_;
  assign new_n485_ = keyinput29 & ~new_n484_;
  assign new_n486_ = ~keyinput29 & new_n484_;
  assign new_n487_ = ~new_n485_ & ~new_n486_;
  assign new_n488_ = ~G4 & G6;
  assign new_n489_ = ~G5 & ~new_n488_;
  assign new_n490_ = ~G1 & G2;
  assign new_n491_ = keyinput45 & new_n490_;
  assign new_n492_ = ~keyinput45 & ~new_n490_;
  assign new_n493_ = ~new_n491_ & ~new_n492_;
  assign new_n494_ = ~new_n489_ & ~new_n493_;
  assign new_n495_ = keyinput25 & ~new_n494_;
  assign new_n496_ = ~keyinput25 & new_n494_;
  assign new_n497_ = ~new_n495_ & ~new_n496_;
  assign new_n498_ = ~new_n478_ & ~new_n487_;
  assign new_n499_ = ~new_n497_ & new_n498_;
  assign new_n500_ = keyinput46 & ~new_n499_;
  assign new_n501_ = ~keyinput46 & new_n499_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = ~new_n296_ & ~new_n502_;
  assign new_n504_ = keyinput75 & ~new_n503_;
  assign new_n505_ = ~keyinput75 & new_n503_;
  assign new_n506_ = ~new_n504_ & ~new_n505_;
  assign new_n507_ = ~G12 & G13;
  assign new_n508_ = new_n506_ & new_n507_;
  assign new_n509_ = new_n460_ & new_n508_;
  assign new_n510_ = new_n312_ & new_n420_;
  assign G539 = new_n509_ | ~new_n510_;
  assign new_n512_ = G5 & ~new_n482_;
  assign new_n513_ = new_n503_ & new_n512_;
  assign new_n514_ = keyinput61 & ~new_n513_;
  assign new_n515_ = ~keyinput61 & new_n513_;
  assign new_n516_ = ~new_n514_ & ~new_n515_;
  assign new_n517_ = new_n482_ & new_n503_;
  assign new_n518_ = ~G5 & new_n517_;
  assign new_n519_ = ~new_n516_ & ~new_n518_;
  assign new_n520_ = G2 & ~new_n519_;
  assign new_n521_ = new_n507_ & new_n520_;
  assign new_n522_ = G2 & G4;
  assign new_n523_ = ~G12 & new_n303_;
  assign new_n524_ = ~G13 & new_n523_;
  assign new_n525_ = keyinput67 & new_n524_;
  assign new_n526_ = ~keyinput67 & ~new_n524_;
  assign new_n527_ = ~new_n525_ & ~new_n526_;
  assign new_n528_ = new_n243_ & ~new_n522_;
  assign new_n529_ = ~new_n527_ & new_n528_;
  assign new_n530_ = keyinput8 & new_n529_;
  assign new_n531_ = ~keyinput8 & ~new_n529_;
  assign new_n532_ = ~new_n530_ & ~new_n531_;
  assign new_n533_ = ~G0 & new_n482_;
  assign new_n534_ = G3 & new_n533_;
  assign new_n535_ = G0 & ~G29;
  assign new_n536_ = ~new_n534_ & ~new_n535_;
  assign new_n537_ = G12 & new_n411_;
  assign new_n538_ = ~G13 & new_n537_;
  assign new_n539_ = keyinput17 & ~new_n538_;
  assign new_n540_ = ~keyinput17 & new_n538_;
  assign new_n541_ = ~new_n539_ & ~new_n540_;
  assign new_n542_ = ~new_n536_ & ~new_n541_;
  assign new_n543_ = keyinput89 & ~G33;
  assign new_n544_ = ~keyinput89 & G33;
  assign new_n545_ = ~new_n543_ & ~new_n544_;
  assign new_n546_ = G3 & ~G13;
  assign new_n547_ = ~new_n545_ & new_n546_;
  assign new_n548_ = keyinput101 & ~new_n547_;
  assign new_n549_ = ~keyinput101 & new_n547_;
  assign new_n550_ = ~new_n548_ & ~new_n549_;
  assign new_n551_ = keyinput85 & new_n550_;
  assign new_n552_ = ~keyinput85 & ~new_n550_;
  assign new_n553_ = ~new_n551_ & ~new_n552_;
  assign new_n554_ = ~new_n521_ & new_n532_;
  assign new_n555_ = ~new_n542_ & new_n554_;
  assign new_n556_ = new_n553_ & new_n555_;
  assign new_n557_ = keyinput21 & ~new_n556_;
  assign new_n558_ = ~keyinput21 & new_n556_;
  assign G550 = new_n557_ | new_n558_;
  assign new_n560_ = G4 & G39;
  assign new_n561_ = ~new_n527_ & new_n560_;
  assign new_n562_ = G0 & G3;
  assign new_n563_ = keyinput18 & new_n562_;
  assign new_n564_ = ~keyinput18 & ~new_n562_;
  assign new_n565_ = ~new_n563_ & ~new_n564_;
  assign new_n566_ = ~new_n482_ & new_n565_;
  assign new_n567_ = G0 & G2;
  assign new_n568_ = G1 & ~new_n567_;
  assign new_n569_ = G4 & new_n567_;
  assign new_n570_ = ~new_n568_ & ~new_n569_;
  assign new_n571_ = ~G3 & ~new_n570_;
  assign new_n572_ = ~new_n566_ & ~new_n571_;
  assign new_n573_ = ~new_n533_ & new_n572_;
  assign new_n574_ = keyinput2 & new_n573_;
  assign new_n575_ = ~keyinput2 & ~new_n573_;
  assign new_n576_ = ~new_n574_ & ~new_n575_;
  assign new_n577_ = G5 & ~new_n576_;
  assign new_n578_ = ~new_n541_ & new_n577_;
  assign new_n579_ = ~G1 & new_n522_;
  assign new_n580_ = new_n503_ & new_n579_;
  assign new_n581_ = keyinput66 & ~new_n517_;
  assign new_n582_ = ~keyinput66 & new_n517_;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign new_n584_ = new_n465_ & new_n583_;
  assign new_n585_ = ~new_n580_ & ~new_n584_;
  assign new_n586_ = keyinput86 & ~new_n585_;
  assign new_n587_ = ~keyinput86 & new_n585_;
  assign new_n588_ = ~new_n586_ & ~new_n587_;
  assign new_n589_ = G6 & new_n465_;
  assign new_n590_ = ~G5 & new_n589_;
  assign new_n591_ = ~G3 & new_n234_;
  assign new_n592_ = ~new_n397_ & ~new_n590_;
  assign new_n593_ = ~new_n591_ & new_n592_;
  assign new_n594_ = G1 & new_n503_;
  assign new_n595_ = ~new_n593_ & new_n594_;
  assign new_n596_ = new_n588_ & ~new_n595_;
  assign new_n597_ = keyinput15 & new_n596_;
  assign new_n598_ = ~keyinput15 & ~new_n596_;
  assign new_n599_ = ~new_n597_ & ~new_n598_;
  assign new_n600_ = new_n507_ & ~new_n599_;
  assign new_n601_ = ~new_n561_ & ~new_n578_;
  assign G551 = new_n600_ | ~new_n601_;
  assign new_n603_ = G2 & G5;
  assign new_n604_ = new_n234_ & ~new_n603_;
  assign new_n605_ = G4 & keyinput71;
  assign new_n606_ = ~G4 & ~keyinput71;
  assign new_n607_ = ~new_n605_ & ~new_n606_;
  assign new_n608_ = G1 & new_n607_;
  assign new_n609_ = G2 & ~new_n608_;
  assign new_n610_ = ~new_n243_ & ~new_n609_;
  assign new_n611_ = G6 & ~new_n610_;
  assign new_n612_ = ~new_n604_ & ~new_n611_;
  assign new_n613_ = ~new_n506_ & ~new_n612_;
  assign new_n614_ = new_n507_ & new_n613_;
  assign new_n615_ = keyinput1 & ~G40;
  assign new_n616_ = ~keyinput1 & G40;
  assign new_n617_ = ~new_n615_ & ~new_n616_;
  assign new_n618_ = ~new_n541_ & new_n617_;
  assign new_n619_ = ~new_n397_ & new_n589_;
  assign new_n620_ = ~G4 & G5;
  assign new_n621_ = ~new_n397_ & ~new_n620_;
  assign new_n622_ = keyinput24 & ~new_n621_;
  assign new_n623_ = ~keyinput24 & new_n621_;
  assign new_n624_ = ~new_n622_ & ~new_n623_;
  assign new_n625_ = G6 & new_n624_;
  assign new_n626_ = ~new_n591_ & ~new_n625_;
  assign new_n627_ = G2 & ~new_n626_;
  assign new_n628_ = keyinput59 & new_n627_;
  assign new_n629_ = ~keyinput59 & ~new_n627_;
  assign new_n630_ = ~new_n628_ & ~new_n629_;
  assign new_n631_ = ~new_n619_ & new_n630_;
  assign new_n632_ = ~new_n527_ & ~new_n631_;
  assign new_n633_ = ~new_n614_ & ~new_n618_;
  assign G552 = new_n632_ | ~new_n633_;
  assign new_n635_ = ~G7 & new_n367_;
  assign new_n636_ = G7 & ~new_n367_;
  assign new_n637_ = keyinput123 & ~new_n636_;
  assign new_n638_ = ~keyinput123 & new_n636_;
  assign new_n639_ = ~new_n637_ & ~new_n638_;
  assign new_n640_ = ~new_n635_ & ~new_n639_;
  assign new_n641_ = keyinput51 & ~G34;
  assign new_n642_ = ~keyinput51 & G34;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign new_n644_ = G9 & ~new_n640_;
  assign new_n645_ = ~new_n643_ & new_n644_;
  assign new_n646_ = ~G6 & new_n249_;
  assign new_n647_ = G9 & new_n646_;
  assign new_n648_ = ~G8 & ~new_n247_;
  assign new_n649_ = G9 & new_n217_;
  assign new_n650_ = ~G10 & new_n233_;
  assign new_n651_ = keyinput40 & ~new_n650_;
  assign new_n652_ = ~keyinput40 & new_n650_;
  assign new_n653_ = ~new_n651_ & ~new_n652_;
  assign new_n654_ = ~new_n649_ & ~new_n653_;
  assign new_n655_ = ~new_n214_ & ~new_n654_;
  assign new_n656_ = ~new_n211_ & new_n218_;
  assign new_n657_ = ~new_n648_ & ~new_n655_;
  assign new_n658_ = ~new_n656_ & new_n657_;
  assign new_n659_ = keyinput6 & ~new_n658_;
  assign new_n660_ = ~keyinput6 & new_n658_;
  assign new_n661_ = ~new_n659_ & ~new_n660_;
  assign new_n662_ = G6 & ~new_n661_;
  assign new_n663_ = ~new_n647_ & ~new_n662_;
  assign new_n664_ = ~new_n541_ & ~new_n663_;
  assign G547 = new_n645_ | new_n664_;
  assign new_n666_ = keyinput58 & ~G42;
  assign new_n667_ = ~keyinput58 & G42;
  assign new_n668_ = ~new_n666_ & ~new_n667_;
  assign new_n669_ = ~new_n541_ & new_n668_;
  assign new_n670_ = new_n244_ & new_n639_;
  assign new_n671_ = ~G9 & new_n249_;
  assign new_n672_ = new_n211_ & ~new_n218_;
  assign new_n673_ = keyinput78 & new_n672_;
  assign new_n674_ = ~keyinput78 & ~new_n672_;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign new_n676_ = ~new_n671_ & ~new_n675_;
  assign new_n677_ = G11 & ~new_n676_;
  assign new_n678_ = ~new_n670_ & ~new_n677_;
  assign new_n679_ = keyinput60 & new_n678_;
  assign new_n680_ = ~keyinput60 & ~new_n678_;
  assign new_n681_ = ~new_n679_ & ~new_n680_;
  assign new_n682_ = ~new_n643_ & ~new_n681_;
  assign G548 = new_n669_ | new_n682_;
  assign new_n684_ = new_n482_ & ~new_n565_;
  assign new_n685_ = ~new_n541_ & new_n684_;
  assign new_n686_ = keyinput43 & ~new_n685_;
  assign new_n687_ = ~keyinput43 & new_n685_;
  assign new_n688_ = ~new_n686_ & ~new_n687_;
  assign new_n689_ = G3 & G4;
  assign new_n690_ = new_n603_ & ~new_n689_;
  assign new_n691_ = ~new_n527_ & new_n690_;
  assign new_n692_ = ~new_n465_ & ~new_n591_;
  assign new_n693_ = G5 & ~new_n692_;
  assign new_n694_ = G2 & new_n397_;
  assign new_n695_ = keyinput38 & ~new_n694_;
  assign new_n696_ = ~keyinput38 & new_n694_;
  assign new_n697_ = ~new_n695_ & ~new_n696_;
  assign new_n698_ = ~G5 & keyinput77;
  assign new_n699_ = G5 & ~keyinput77;
  assign new_n700_ = ~new_n698_ & ~new_n699_;
  assign new_n701_ = ~new_n466_ & ~new_n700_;
  assign new_n702_ = ~G4 & ~new_n701_;
  assign new_n703_ = ~new_n693_ & ~new_n697_;
  assign new_n704_ = ~new_n702_ & new_n703_;
  assign new_n705_ = new_n507_ & ~new_n704_;
  assign new_n706_ = new_n594_ & new_n705_;
  assign new_n707_ = keyinput70 & ~new_n706_;
  assign new_n708_ = ~keyinput70 & new_n706_;
  assign new_n709_ = ~new_n707_ & ~new_n708_;
  assign new_n710_ = new_n688_ & ~new_n691_;
  assign new_n711_ = new_n709_ & new_n710_;
  assign G549 = new_n550_ | ~new_n711_;
  assign new_n713_ = ~G0 & G1;
  assign new_n714_ = ~G5 & new_n421_;
  assign new_n715_ = ~G4 & new_n243_;
  assign new_n716_ = ~new_n714_ & ~new_n715_;
  assign new_n717_ = ~new_n389_1_ & new_n716_;
  assign new_n718_ = keyinput93 & ~new_n717_;
  assign new_n719_ = ~keyinput93 & new_n717_;
  assign new_n720_ = ~new_n718_ & ~new_n719_;
  assign new_n721_ = G0 & ~new_n720_;
  assign new_n722_ = ~new_n713_ & ~new_n721_;
  assign new_n723_ = keyinput33 & ~new_n722_;
  assign new_n724_ = ~keyinput33 & new_n722_;
  assign new_n725_ = ~new_n723_ & ~new_n724_;
  assign new_n726_ = G2 & ~new_n725_;
  assign new_n727_ = ~new_n541_ & new_n726_;
  assign new_n728_ = ~new_n291_ & new_n307_;
  assign new_n729_ = ~G12 & new_n728_;
  assign new_n730_ = ~new_n288_ & new_n729_;
  assign new_n731_ = keyinput65 & new_n730_;
  assign new_n732_ = ~keyinput65 & ~new_n730_;
  assign new_n733_ = ~new_n731_ & ~new_n732_;
  assign G530 = new_n727_ | ~new_n733_;
  assign new_n735_ = G8 & G9;
  assign new_n736_ = new_n249_ & ~new_n735_;
  assign new_n737_ = ~new_n643_ & new_n736_;
  assign new_n738_ = G7 & G9;
  assign new_n739_ = keyinput90 & ~new_n738_;
  assign new_n740_ = ~keyinput90 & new_n738_;
  assign new_n741_ = ~new_n739_ & ~new_n740_;
  assign new_n742_ = new_n367_ & ~new_n741_;
  assign new_n743_ = keyinput28 & new_n742_;
  assign new_n744_ = ~keyinput28 & ~new_n742_;
  assign new_n745_ = ~new_n743_ & ~new_n744_;
  assign new_n746_ = G7 & ~G8;
  assign new_n747_ = keyinput69 & ~new_n746_;
  assign new_n748_ = ~keyinput69 & new_n746_;
  assign new_n749_ = ~new_n747_ & ~new_n748_;
  assign new_n750_ = keyinput32 & ~new_n217_;
  assign new_n751_ = ~keyinput32 & new_n217_;
  assign new_n752_ = ~new_n750_ & ~new_n751_;
  assign new_n753_ = keyinput76 & ~new_n752_;
  assign new_n754_ = ~keyinput76 & new_n752_;
  assign new_n755_ = ~new_n753_ & ~new_n754_;
  assign new_n756_ = ~new_n749_ & ~new_n755_;
  assign new_n757_ = ~G9 & ~new_n756_;
  assign new_n758_ = ~new_n429_ & ~new_n745_;
  assign new_n759_ = ~new_n757_ & new_n758_;
  assign new_n760_ = keyinput119 & ~new_n759_;
  assign new_n761_ = ~keyinput119 & new_n759_;
  assign new_n762_ = ~new_n760_ & ~new_n761_;
  assign new_n763_ = G6 & ~new_n541_;
  assign new_n764_ = new_n762_ & new_n763_;
  assign new_n765_ = G8 & ~new_n643_;
  assign new_n766_ = ~new_n763_ & ~new_n765_;
  assign new_n767_ = new_n294_ & ~new_n766_;
  assign new_n768_ = ~new_n737_ & ~new_n764_;
  assign G542 = new_n767_ | ~new_n768_;
  assign new_n770_ = ~G3 & keyinput114;
  assign new_n771_ = G3 & ~keyinput114;
  assign new_n772_ = ~new_n770_ & ~new_n771_;
  assign new_n773_ = G1 & ~G2;
  assign new_n774_ = new_n772_ & new_n773_;
  assign new_n775_ = ~G3 & ~G5;
  assign new_n776_ = G2 & ~new_n421_;
  assign new_n777_ = ~G2 & new_n243_;
  assign new_n778_ = keyinput124 & ~new_n777_;
  assign new_n779_ = ~keyinput124 & new_n777_;
  assign new_n780_ = ~new_n778_ & ~new_n779_;
  assign new_n781_ = ~new_n775_ & ~new_n776_;
  assign new_n782_ = ~new_n780_ & new_n781_;
  assign new_n783_ = G4 & ~new_n782_;
  assign new_n784_ = ~new_n422_ & ~new_n774_;
  assign new_n785_ = ~new_n783_ & new_n784_;
  assign new_n786_ = G0 & ~new_n785_;
  assign new_n787_ = ~new_n541_ & new_n786_;
  assign new_n788_ = keyinput73 & ~new_n460_;
  assign new_n789_ = ~keyinput73 & new_n460_;
  assign new_n790_ = ~new_n788_ & ~new_n789_;
  assign new_n791_ = G13 & new_n790_;
  assign new_n792_ = keyinput126 & new_n791_;
  assign new_n793_ = ~keyinput126 & ~new_n791_;
  assign new_n794_ = ~new_n792_ & ~new_n793_;
  assign new_n795_ = keyinput63 & new_n794_;
  assign new_n796_ = ~keyinput63 & ~new_n794_;
  assign new_n797_ = ~new_n795_ & ~new_n796_;
  assign new_n798_ = keyinput117 & new_n728_;
  assign new_n799_ = ~keyinput117 & ~new_n728_;
  assign new_n800_ = ~new_n798_ & ~new_n799_;
  assign new_n801_ = new_n797_ & new_n800_;
  assign new_n802_ = ~G4 & ~new_n229_;
  assign new_n803_ = keyinput92 & new_n802_;
  assign new_n804_ = ~keyinput92 & ~new_n802_;
  assign new_n805_ = ~new_n803_ & ~new_n804_;
  assign new_n806_ = keyinput52 & new_n266_;
  assign new_n807_ = ~keyinput52 & ~new_n266_;
  assign new_n808_ = ~new_n806_ & ~new_n807_;
  assign new_n809_ = new_n805_ & ~new_n808_;
  assign new_n810_ = G6 & keyinput37;
  assign new_n811_ = ~G6 & ~keyinput37;
  assign new_n812_ = ~new_n810_ & ~new_n811_;
  assign new_n813_ = ~new_n801_ & ~new_n809_;
  assign new_n814_ = ~new_n812_ & new_n813_;
  assign new_n815_ = keyinput80 & ~new_n794_;
  assign new_n816_ = ~keyinput80 & new_n794_;
  assign new_n817_ = ~new_n815_ & ~new_n816_;
  assign new_n818_ = new_n235_ & new_n728_;
  assign new_n819_ = new_n817_ & ~new_n818_;
  assign new_n820_ = ~new_n432_ & ~new_n819_;
  assign new_n821_ = keyinput35 & ~G43;
  assign new_n822_ = ~keyinput35 & G43;
  assign new_n823_ = ~new_n821_ & ~new_n822_;
  assign new_n824_ = G13 & ~new_n506_;
  assign new_n825_ = new_n823_ & new_n824_;
  assign new_n826_ = keyinput88 & ~new_n825_;
  assign new_n827_ = ~keyinput88 & new_n825_;
  assign new_n828_ = ~new_n826_ & ~new_n827_;
  assign new_n829_ = ~new_n281_ & new_n447_;
  assign new_n830_ = ~new_n441_ & ~new_n829_;
  assign new_n831_ = ~G3 & ~new_n830_;
  assign new_n832_ = new_n728_ & new_n831_;
  assign new_n833_ = ~new_n814_ & ~new_n820_;
  assign new_n834_ = new_n828_ & new_n833_;
  assign new_n835_ = ~new_n832_ & new_n834_;
  assign new_n836_ = ~G12 & ~new_n835_;
  assign G532 = new_n787_ | new_n836_;
  assign new_n838_ = new_n340_ & ~new_n416_;
  assign new_n839_ = new_n454_ & new_n838_;
  assign new_n840_ = G37 & new_n839_;
  assign new_n841_ = G38 & new_n840_;
  assign new_n842_ = keyinput79 & ~new_n218_;
  assign new_n843_ = ~keyinput79 & new_n218_;
  assign new_n844_ = ~new_n842_ & ~new_n843_;
  assign new_n845_ = ~new_n227_ & ~new_n844_;
  assign new_n846_ = new_n397_ & ~new_n817_;
  assign new_n847_ = ~new_n845_ & new_n846_;
  assign new_n848_ = ~new_n801_ & ~new_n805_;
  assign new_n849_ = ~new_n847_ & ~new_n848_;
  assign new_n850_ = ~G12 & ~new_n849_;
  assign new_n851_ = ~new_n812_ & new_n850_;
  assign new_n852_ = ~new_n841_ & ~new_n851_;
  assign new_n853_ = keyinput9 & new_n852_;
  assign new_n854_ = ~keyinput9 & ~new_n852_;
  assign new_n855_ = ~new_n853_ & ~new_n854_;
  assign new_n856_ = ~new_n240_ & ~new_n845_;
  assign new_n857_ = keyinput110 & ~G44;
  assign new_n858_ = ~keyinput110 & G44;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = ~G3 & new_n859_;
  assign new_n861_ = ~new_n856_ & ~new_n860_;
  assign new_n862_ = keyinput125 & ~new_n861_;
  assign new_n863_ = ~keyinput125 & new_n861_;
  assign new_n864_ = ~new_n862_ & ~new_n863_;
  assign new_n865_ = new_n729_ & ~new_n864_;
  assign G535 = new_n855_ | new_n865_;
  assign new_n867_ = new_n227_ & ~new_n812_;
  assign new_n868_ = keyinput104 & ~new_n867_;
  assign new_n869_ = ~keyinput104 & new_n867_;
  assign new_n870_ = ~new_n868_ & ~new_n869_;
  assign new_n871_ = keyinput62 & new_n243_;
  assign new_n872_ = ~keyinput62 & ~new_n243_;
  assign new_n873_ = ~new_n871_ & ~new_n872_;
  assign new_n874_ = new_n870_ & new_n873_;
  assign new_n875_ = G8 & ~new_n801_;
  assign new_n876_ = ~new_n874_ & new_n875_;
  assign new_n877_ = keyinput122 & new_n876_;
  assign new_n878_ = ~keyinput122 & ~new_n876_;
  assign new_n879_ = ~new_n877_ & ~new_n878_;
  assign new_n880_ = keyinput3 & new_n229_;
  assign new_n881_ = ~keyinput3 & ~new_n229_;
  assign new_n882_ = ~new_n880_ & ~new_n881_;
  assign new_n883_ = new_n235_ & new_n882_;
  assign new_n884_ = ~new_n817_ & new_n883_;
  assign new_n885_ = keyinput26 & ~new_n884_;
  assign new_n886_ = ~keyinput26 & new_n884_;
  assign new_n887_ = ~new_n885_ & ~new_n886_;
  assign new_n888_ = new_n879_ & new_n887_;
  assign new_n889_ = keyinput98 & ~new_n888_;
  assign new_n890_ = ~keyinput98 & new_n888_;
  assign new_n891_ = ~new_n889_ & ~new_n890_;
  assign new_n892_ = ~G12 & ~new_n891_;
  assign new_n893_ = G38 & new_n317_;
  assign new_n894_ = ~new_n249_ & ~new_n893_;
  assign new_n895_ = keyinput108 & ~new_n894_;
  assign new_n896_ = ~keyinput108 & new_n894_;
  assign new_n897_ = ~new_n895_ & ~new_n896_;
  assign new_n898_ = new_n839_ & ~new_n897_;
  assign new_n899_ = ~new_n892_ & ~new_n898_;
  assign new_n900_ = G2 & ~new_n899_;
  assign new_n901_ = keyinput30 & new_n900_;
  assign new_n902_ = ~keyinput30 & ~new_n900_;
  assign new_n903_ = ~new_n901_ & ~new_n902_;
  assign new_n904_ = new_n248_ & new_n397_;
  assign new_n905_ = new_n646_ & new_n904_;
  assign new_n906_ = ~G5 & new_n441_;
  assign new_n907_ = new_n344_1_ & new_n906_;
  assign new_n908_ = G10 & ~new_n247_;
  assign new_n909_ = ~new_n281_ & new_n908_;
  assign new_n910_ = ~new_n907_ & ~new_n909_;
  assign new_n911_ = ~new_n378_ & ~new_n910_;
  assign new_n912_ = keyinput100 & new_n911_;
  assign new_n913_ = ~keyinput100 & ~new_n911_;
  assign new_n914_ = ~new_n912_ & ~new_n913_;
  assign new_n915_ = ~new_n905_ & new_n914_;
  assign new_n916_ = ~new_n883_ & new_n915_;
  assign new_n917_ = new_n729_ & ~new_n916_;
  assign new_n918_ = keyinput74 & new_n917_;
  assign new_n919_ = ~keyinput74 & ~new_n917_;
  assign new_n920_ = ~new_n918_ & ~new_n919_;
  assign new_n921_ = new_n903_ & new_n920_;
  assign new_n922_ = keyinput31 & new_n921_;
  assign new_n923_ = ~keyinput31 & ~new_n921_;
  assign G537 = new_n922_ | new_n923_;
  assign new_n925_ = ~new_n397_ & new_n465_;
  assign new_n926_ = keyinput42 & new_n925_;
  assign new_n927_ = ~keyinput42 & ~new_n925_;
  assign new_n928_ = ~new_n926_ & ~new_n927_;
  assign new_n929_ = ~new_n620_ & ~new_n689_;
  assign new_n930_ = ~new_n493_ & ~new_n929_;
  assign n314 = new_n928_ & ~new_n930_;
  assign new_n932_ = ~G9 & new_n233_;
  assign n319 = new_n217_ | new_n932_;
  assign new_n934_ = new_n217_ & new_n247_;
  assign new_n935_ = keyinput64 & ~new_n934_;
  assign new_n936_ = ~keyinput64 & new_n934_;
  assign new_n937_ = ~new_n935_ & ~new_n936_;
  assign new_n938_ = ~G7 & new_n233_;
  assign new_n939_ = ~new_n937_ & ~new_n938_;
  assign new_n940_ = keyinput44 & new_n939_;
  assign new_n941_ = ~keyinput44 & ~new_n939_;
  assign n324 = new_n940_ | new_n941_;
  assign new_n943_ = ~new_n235_ & new_n603_;
  assign new_n944_ = keyinput20 & ~new_n943_;
  assign new_n945_ = ~keyinput20 & new_n943_;
  assign new_n946_ = ~new_n944_ & ~new_n945_;
  assign new_n947_ = new_n465_ & ~new_n489_;
  assign new_n948_ = ~new_n946_ & ~new_n947_;
  assign n329 = new_n697_ | ~new_n948_;
  assign new_n950_ = G1 & ~G4;
  assign new_n951_ = G0 & new_n950_;
  assign new_n952_ = new_n537_ & new_n951_;
  assign new_n953_ = new_n523_ & new_n697_;
  assign n334 = ~new_n952_ & ~new_n953_;
  assign new_n955_ = G13 & ~new_n502_;
  assign new_n956_ = ~G13 & ~new_n299_;
  assign new_n957_ = ~new_n955_ & ~new_n956_;
  assign new_n958_ = ~G12 & ~new_n957_;
  assign n339 = ~new_n296_ & new_n958_;
  assign new_n960_ = ~G6 & ~G8;
  assign new_n961_ = new_n227_ & new_n960_;
  assign new_n962_ = keyinput10 & ~new_n961_;
  assign new_n963_ = ~keyinput10 & new_n961_;
  assign new_n964_ = ~new_n962_ & ~new_n963_;
  assign new_n965_ = G6 & ~new_n229_;
  assign n344 = new_n964_ | new_n965_;
  assign new_n967_ = ~new_n217_ & ~new_n264_;
  assign new_n968_ = keyinput11 & new_n967_;
  assign new_n969_ = ~keyinput11 & ~new_n967_;
  assign new_n970_ = ~new_n968_ & ~new_n969_;
  assign new_n971_ = ~new_n250_ & ~new_n970_;
  assign new_n972_ = ~G5 & ~new_n971_;
  assign new_n973_ = keyinput107 & ~new_n972_;
  assign new_n974_ = ~keyinput107 & new_n972_;
  assign n349 = new_n973_ | new_n974_;
  assign new_n976_ = ~G6 & G9;
  assign n354 = new_n317_ | new_n976_;
  assign n359 = new_n226_ & new_n328_;
  assign new_n979_ = G2 & ~new_n243_;
  assign n364 = new_n780_ | new_n979_;
  assign new_n981_ = G6 & G9;
  assign new_n982_ = ~G11 & new_n981_;
  assign new_n983_ = ~G6 & G30;
  assign new_n984_ = ~new_n982_ & ~new_n983_;
  assign new_n985_ = G7 & ~new_n984_;
  assign new_n986_ = keyinput87 & ~new_n985_;
  assign new_n987_ = ~keyinput87 & new_n985_;
  assign new_n988_ = ~new_n986_ & ~new_n987_;
  assign new_n989_ = G6 & G31;
  assign new_n990_ = new_n988_ & ~new_n989_;
  assign new_n991_ = G8 & ~new_n990_;
  assign new_n992_ = G6 & ~new_n437_;
  assign n369 = ~new_n991_ & ~new_n992_;
  assign new_n994_ = new_n249_ & ~new_n981_;
  assign new_n995_ = ~new_n541_ & new_n994_;
  assign new_n996_ = keyinput102 & ~new_n745_;
  assign new_n997_ = ~keyinput102 & new_n745_;
  assign new_n998_ = ~new_n996_ & ~new_n997_;
  assign new_n999_ = ~new_n643_ & ~new_n998_;
  assign new_n1000_ = keyinput72 & new_n999_;
  assign new_n1001_ = ~keyinput72 & ~new_n999_;
  assign new_n1002_ = ~new_n1000_ & ~new_n1001_;
  assign new_n1003_ = ~new_n995_ & new_n1002_;
  assign n374 = ~new_n767_ & new_n1003_;
  assign new_n1005_ = G6 & ~new_n249_;
  assign new_n1006_ = ~new_n247_ & new_n1005_;
  assign new_n1007_ = ~new_n218_ & new_n349_1_;
  assign new_n1008_ = G6 & new_n367_;
  assign new_n1009_ = keyinput39 & new_n1008_;
  assign new_n1010_ = ~keyinput39 & ~new_n1008_;
  assign new_n1011_ = ~new_n1009_ & ~new_n1010_;
  assign new_n1012_ = ~new_n749_ & ~new_n1011_;
  assign new_n1013_ = ~G9 & ~new_n1012_;
  assign new_n1014_ = ~new_n1007_ & ~new_n1013_;
  assign new_n1015_ = G11 & ~new_n1014_;
  assign n379 = ~new_n1006_ & ~new_n1015_;
  assign new_n1017_ = G1 & new_n589_;
  assign new_n1018_ = ~G6 & new_n522_;
  assign new_n1019_ = G6 & new_n397_;
  assign new_n1020_ = keyinput84 & ~new_n1019_;
  assign new_n1021_ = ~keyinput84 & new_n1019_;
  assign new_n1022_ = ~new_n1020_ & ~new_n1021_;
  assign new_n1023_ = G5 & ~new_n234_;
  assign new_n1024_ = ~new_n1018_ & ~new_n1022_;
  assign new_n1025_ = ~new_n1023_ & new_n1024_;
  assign new_n1026_ = keyinput41 & ~new_n1025_;
  assign new_n1027_ = ~keyinput41 & new_n1025_;
  assign new_n1028_ = ~new_n1026_ & ~new_n1027_;
  assign new_n1029_ = new_n421_ & ~new_n1028_;
  assign new_n1030_ = keyinput116 & ~new_n1029_;
  assign new_n1031_ = ~keyinput116 & new_n1029_;
  assign new_n1032_ = ~new_n1030_ & ~new_n1031_;
  assign new_n1033_ = G3 & new_n497_;
  assign new_n1034_ = ~new_n1017_ & new_n1032_;
  assign n384 = ~new_n1033_ & new_n1034_;
  assign new_n1036_ = new_n250_ & new_n906_;
  assign new_n1037_ = ~G5 & ~G6;
  assign new_n1038_ = new_n348_ & new_n1037_;
  assign new_n1039_ = ~new_n909_ & ~new_n1038_;
  assign new_n1040_ = ~new_n378_ & ~new_n1039_;
  assign n389 = ~new_n1036_ & ~new_n1040_;
  assign new_n1042_ = ~new_n460_ & new_n508_;
  assign new_n1043_ = keyinput94 & ~new_n1042_;
  assign new_n1044_ = ~keyinput94 & new_n1042_;
  assign new_n1045_ = ~new_n1043_ & ~new_n1044_;
  assign new_n1046_ = ~new_n729_ & ~new_n838_;
  assign n394 = new_n1045_ | ~new_n1046_;
  assign new_n1048_ = G0 & G4;
  assign new_n1049_ = keyinput106 & new_n442_;
  assign new_n1050_ = ~keyinput106 & ~new_n442_;
  assign new_n1051_ = ~new_n1049_ & ~new_n1050_;
  assign new_n1052_ = keyinput14 & new_n1051_;
  assign new_n1053_ = ~keyinput14 & ~new_n1051_;
  assign new_n1054_ = ~new_n1052_ & ~new_n1053_;
  assign new_n1055_ = G0 & ~G3;
  assign new_n1056_ = ~new_n1048_ & new_n1054_;
  assign new_n1057_ = ~new_n1055_ & new_n1056_;
  assign new_n1058_ = G2 & ~new_n389_1_;
  assign new_n1059_ = ~new_n1057_ & new_n1058_;
  assign new_n1060_ = ~G6 & ~G7;
  assign new_n1061_ = keyinput36 & new_n1060_;
  assign new_n1062_ = ~keyinput36 & ~new_n1060_;
  assign new_n1063_ = ~new_n1061_ & ~new_n1062_;
  assign new_n1064_ = ~new_n217_ & new_n374_1_;
  assign new_n1065_ = new_n397_ & new_n465_;
  assign new_n1066_ = new_n391_ & ~new_n397_;
  assign new_n1067_ = ~new_n1065_ & ~new_n1066_;
  assign new_n1068_ = G0 & new_n1067_;
  assign new_n1069_ = ~G1 & ~new_n1068_;
  assign new_n1070_ = ~new_n1059_ & new_n1063_;
  assign new_n1071_ = ~new_n1064_ & new_n1070_;
  assign n398 = ~new_n1069_ & new_n1071_;
  assign G546 = ~G41;
  always @ (posedge clock) begin
    G29 <= n314;
    G30 <= n319;
    G31 <= n324;
    G32 <= n329;
    G33 <= n334;
    G34 <= n339;
    G35 <= n344;
    G36 <= n349;
    G37 <= n354;
    G38 <= n359;
    G39 <= n364;
    G40 <= n369;
    G41 <= n374;
    G42 <= n379;
    G43 <= n384;
    G44 <= n389;
    G45 <= n394;
    G46 <= n398;
  end
endmodule


